/**
 * eth.sv:
 *   This file wraps Ethernet controller module with AXI
 */

module eth #(
    parameter burst_size = 16,
    parameter dma_word_bits = 32,
    parameter dma_addr_bits = 32,
    parameter axis_word_bits = 8,
    parameter pkt_ptr_bits = 4, /* max is 6 */
    parameter enable_mdio = 1,
    parameter blk = 64 // cache block size
)(
    input  logic        clk,
    input  logic        rst,
    input  logic [15:0] status_vector,
    output logic        intr,
    output logic        rst_o,
    /* AXI slave interface */
    input  logic [15:0] s_axi_awaddr,
    input  logic        s_axi_awvalid,
    output logic        s_axi_awready,
    input  logic [31:0] s_axi_wdata,
    input  logic        s_axi_wvalid,
    output logic        s_axi_wready,
    output logic  [1:0] s_axi_bresp,
    output logic        s_axi_bvalid,
    input  logic        s_axi_bready,
    input  logic [15:0] s_axi_araddr,
    input  logic        s_axi_arvalid,
    output logic        s_axi_arready,
    output logic [31:0] s_axi_rdata,
    output logic  [1:0] s_axi_rresp,
    output logic        s_axi_rvalid,
    input  logic        s_axi_rready,
    /* AXI master interface */
    output logic   [dma_addr_bits-1:0] m_axi_awaddr,
    output logic                 [7:0] m_axi_awlen,
    output logic                 [2:0] m_axi_awsize,
    output logic                 [1:0] m_axi_awburst,
    output logic                       m_axi_awvalid,
    input  logic                       m_axi_awready,
    output logic   [dma_word_bits-1:0] m_axi_wdata,
    output logic [dma_word_bits/8-1:0] m_axi_wstrb,
    output logic                       m_axi_wlast,
    output logic                       m_axi_wvalid,
    input  logic                       m_axi_wready,
    input  logic                 [1:0] m_axi_bresp,
    input  logic                       m_axi_bvalid,
    output logic                       m_axi_bready,
    output logic   [dma_addr_bits-1:0] m_axi_araddr,
    output logic                 [7:0] m_axi_arlen,
    output logic                 [2:0] m_axi_arsize,
    output logic                 [1:0] m_axi_arburst,
    output logic                       m_axi_arvalid,
    input  logic                       m_axi_arready,
    input  logic   [dma_word_bits-1:0] m_axi_rdata,
    input  logic                       m_axi_rlast,
    input  logic                 [1:0] m_axi_rresp,
    input  logic                       m_axi_rvalid,
    output logic                       m_axi_rready,
    /* TX interface */
    output logic   [axis_word_bits-1:0] tx_axis_tdata,
    output logic [axis_word_bits/8-1:0] tx_axis_tkeep,
    output logic                        tx_axis_tvalid,
    input  logic                        tx_axis_tready,
    output logic                        tx_axis_tlast,
    output logic                        tx_axis_tuser,
    /* RX interface */
    input  logic   [axis_word_bits-1:0] rx_axis_tdata,
    input  logic [axis_word_bits/8-1:0] rx_axis_tkeep,
    input  logic                        rx_axis_tvalid,
    output logic                        rx_axis_tready,
    input  logic                        rx_axis_tlast,
    input  logic                        rx_axis_tuser,
    /* MDIO interface */
    output logic mdio_clock,
    output logic mdio_data_t,
    output logic mdio_data_o,
    input  logic mdio_data_i,
    output logic mdio_reset,
    input  logic mdio_int
);
    /* instance */
    ethernet ethernet_inst(
        .clock(clk),
        .async_resetn(~rst),
        .status_vector(status_vector),
        .interrupt(intr),
        .reset(rst_o),
        .s_axi_awaddr(s_axi_awaddr),
        .s_axi_awvalid(s_axi_awvalid),
        .s_axi_awready(s_axi_awready),
        .s_axi_wdata(s_axi_wdata),
        .s_axi_wvalid(s_axi_wvalid),
        .s_axi_wready(s_axi_wready),
        .s_axi_bresp(s_axi_bresp),
        .s_axi_bvalid(s_axi_bvalid),
        .s_axi_bready(s_axi_bready),
        .s_axi_araddr(s_axi_araddr),
        .s_axi_arvalid(s_axi_arvalid),
        .s_axi_arready(s_axi_arready),
        .s_axi_rdata(s_axi_rdata),
        .s_axi_rresp(s_axi_rresp),
        .s_axi_rvalid(s_axi_rvalid),
        .s_axi_rready(s_axi_rready),
        .m_axi_awaddr(m_axi_awaddr),
        .m_axi_awlen(m_axi_awlen),
        .m_axi_awvalid(m_axi_awvalid),
        .m_axi_awready(m_axi_awready),
        .m_axi_wdata(m_axi_wdata),
        .m_axi_wstrb(m_axi_wstrb),
        .m_axi_wlast(m_axi_wlast),
        .m_axi_wvalid(m_axi_wvalid),
        .m_axi_wready(m_axi_wready),
        .m_axi_bresp(m_axi_bresp),
        .m_axi_bvalid(m_axi_bvalid),
        .m_axi_bready(m_axi_bready),
        .m_axi_araddr(m_axi_araddr),
        .m_axi_arlen(m_axi_arlen),
        .m_axi_arvalid(m_axi_arvalid),
        .m_axi_arready(m_axi_arready),
        .m_axi_rdata(m_axi_rdata),
        .m_axi_rlast(m_axi_rlast),
        .m_axi_rresp(m_axi_rresp),
        .m_axi_rvalid(m_axi_rvalid),
        .m_axi_rready(m_axi_rready),
        .tx_axis_tdata(tx_axis_tdata),
        .tx_axis_tkeep(tx_axis_tkeep),
        .tx_axis_tvalid(tx_axis_tvalid),
        .tx_axis_tready(tx_axis_tready),
        .tx_axis_tlast(tx_axis_tlast),
        .tx_axis_tuser(tx_axis_tuser),
        .rx_axis_tdata(rx_axis_tdata),
        .rx_axis_tkeep(rx_axis_tkeep),
        .rx_axis_tvalid(rx_axis_tvalid),
        .rx_axis_tready(rx_axis_tready),
        .rx_axis_tlast(rx_axis_tlast),
        .rx_axis_tuser(rx_axis_tuser),
        .mdio_clock(mdio_clock),
        .mdio_data_t(mdio_data_t),
        .mdio_data_o(mdio_data_o),
        .mdio_data_i(mdio_data_i),
        .mdio_reset(mdio_reset),
        .mdio_int(mdio_int)
    );
    always_comb m_axi_awsize = 2;  // 32-bit
    always_comb m_axi_awburst = 1; // INCR
    always_comb m_axi_arsize = 2;
    always_comb m_axi_arburst = 1;
endmodule
