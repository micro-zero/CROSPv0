/**
 * sdc.sv:
 *   This file wraps SD card controller module with AXI-Lite
 */

module sdc(
    input  logic clk,
    input  logic rst,
    output logic intr,
    /* slave interface for SDC */
    input  logic [15:0] s_axi_awaddr,
    input  logic        s_axi_awvalid,
    output logic        s_axi_awready,
    input  logic [31:0] s_axi_wdata,
    input  logic        s_axi_wvalid,
    output logic        s_axi_wready,
    output logic  [1:0] s_axi_bresp,
    output logic        s_axi_bvalid,
    input  logic        s_axi_bready,
    input  logic [15:0] s_axi_araddr,
    input  logic        s_axi_arvalid,
    output logic        s_axi_arready,
    output logic [31:0] s_axi_rdata,
    output logic  [1:0] s_axi_rresp,
    output logic        s_axi_rvalid,
    input  logic        s_axi_rready,
    /* master interface for SDC */
    output logic [31:0] m_axi_awaddr,
    output logic  [7:0] m_axi_awlen,
    output logic  [2:0] m_axi_awsize,
    output logic  [1:0] m_axi_awburst,
    output logic        m_axi_awvalid,
    input  logic        m_axi_awready,
    output logic [31:0] m_axi_wdata,
    output logic  [3:0] m_axi_wstrb,
    output logic        m_axi_wlast,
    output logic        m_axi_wvalid,
    input  logic        m_axi_wready,
    input  logic  [1:0] m_axi_bresp,
    input  logic        m_axi_bvalid,
    output logic        m_axi_bready,
    output logic [31:0] m_axi_araddr,
    output logic  [7:0] m_axi_arlen,
    output logic  [2:0] m_axi_arsize,
    output logic  [1:0] m_axi_arburst,
    output logic        m_axi_arvalid,
    input  logic        m_axi_arready,
    input  logic [31:0] m_axi_rdata,
    input  logic        m_axi_rlast,
    input  logic  [1:0] m_axi_rresp,
    input  logic        m_axi_rvalid,
    output logic        m_axi_rready,
    /* SD card interface */
    input  logic       sd_cd,
    output logic       sd_cmd_t,
    input  logic       sd_cmd_i,
    output logic       sd_cmd_o,
    output logic       sd_dat_t,
    input  logic [3:0] sd_dat_i,
    output logic [3:0] sd_dat_o,
    output logic       sd_reset,
    output logic       sd_sclk
);
    sdc_controller sdc_inst(
        .clock(clk),
        .async_resetn(~rst),
        .interrupt(intr),
        .s_axi_awaddr(s_axi_awaddr),
        .s_axi_awvalid(s_axi_awvalid),
        .s_axi_awready(s_axi_awready),
        .s_axi_wdata(s_axi_wdata),
        .s_axi_wvalid(s_axi_wvalid),
        .s_axi_wready(s_axi_wready),
        .s_axi_bresp(s_axi_bresp),
        .s_axi_bvalid(s_axi_bvalid),
        .s_axi_bready(s_axi_bready),
        .s_axi_araddr(s_axi_araddr),
        .s_axi_arvalid(s_axi_arvalid),
        .s_axi_arready(s_axi_arready),
        .s_axi_rdata(s_axi_rdata),
        .s_axi_rresp(s_axi_rresp),
        .s_axi_rvalid(s_axi_rvalid),
        .s_axi_rready(s_axi_rready),
        .m_axi_awaddr(m_axi_awaddr),
        .m_axi_awlen(m_axi_awlen),
        .m_axi_awvalid(m_axi_awvalid),
        .m_axi_awready(m_axi_awready),
        .m_axi_wdata(m_axi_wdata),
        .m_axi_wlast(m_axi_wlast),
        .m_axi_wvalid(m_axi_wvalid),
        .m_axi_wready(m_axi_wready),
        .m_axi_bresp(m_axi_bresp),
        .m_axi_bvalid(m_axi_bvalid),
        .m_axi_bready(m_axi_bready),
        .m_axi_araddr(m_axi_araddr),
        .m_axi_arlen(m_axi_arlen),
        .m_axi_arvalid(m_axi_arvalid),
        .m_axi_arready(m_axi_arready),
        .m_axi_rdata(m_axi_rdata),
        .m_axi_rlast(m_axi_rlast),
        .m_axi_rresp(m_axi_rresp),
        .m_axi_rvalid(m_axi_rvalid),
        .m_axi_rready(m_axi_rready),
        .sdio_cd(sd_cd),
        .sd_cmd_reg_t(sd_cmd_t),
        .sd_cmd_i(sd_cmd_i),
        .sd_cmd_reg_o(sd_cmd_o),
        .sd_dat_reg_t(sd_dat_t),
        .sd_dat_i(sd_dat_i),
        .sd_dat_reg_o(sd_dat_o),
        .sdio_reset(sd_reset),
        .sdio_clk(sd_sclk)
    );
    always_comb m_axi_awsize = 2;  // 32-bit
    always_comb m_axi_awburst = 1; // INCR
    always_comb m_axi_arsize = 2;
    always_comb m_axi_arburst = 1;
    always_comb m_axi_wstrb = 'hf;
endmodule
